* C:\Users\vinit\Desktop\SUMMATION-OF-COUNTER\vinit_inverter\vinit_inverter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/21/23 20:28:49

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC2  Net-_SC1-Pad1_ A GND GND sky130_fd_pr__nfet_01v8_lvt		
SC1  Net-_SC1-Pad1_ A Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
v1  Net-_SC1-Pad3_ GND 1.8		
v2  A GND pulse		
scmode1  SKY130mode		
U1  A plot_v1		
U2  y plot_v1		
SC3  Net-_SC1-Pad1_ y Net-_SC1-Pad1_ sky130_fd_pr__res_generic_pd		
SC4  y GND sky130_fd_pr__cap_mim_m3_1		

.end
