* C:\Users\vinit\Desktop\SUMMATION-OF-COUNTER\vinit_2bitpa\vinit_2bitpa.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/29/23 22:48:17

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_U7-Pad1_ GND pulse		
v2  Net-_U7-Pad2_ GND pulse		
v3  Net-_U7-Pad3_ GND pulse		
U11  s1 plot_v1		
U10  s2 plot_v1		
U9  c0 plot_v1		
U7  Net-_U7-Pad1_ Net-_U7-Pad2_ Net-_U7-Pad3_ Net-_U7-Pad4_ GND a1 a2 b1 b2 cin adc_bridge_5		
v4  Net-_U7-Pad4_ GND pulse		
U8  Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_SC3-Pad1_ Net-_SC2-Pad1_ Net-_SC1-Pad1_ dac_bridge_3		
SC3  Net-_SC3-Pad1_ s1 Net-_SC3-Pad1_ sky130_fd_pr__res_generic_pd		
SC2  Net-_SC2-Pad1_ s2 Net-_SC2-Pad1_ sky130_fd_pr__res_generic_pd		
SC1  Net-_SC1-Pad1_ c0 Net-_SC1-Pad1_ sky130_fd_pr__res_generic_pd		
SC6  s1 GND sky130_fd_pr__cap_mim_m3_1		
SC5  s2 GND sky130_fd_pr__cap_mim_m3_1		
SC4  c0 GND sky130_fd_pr__cap_mim_m3_1		
scmode1  SKY130mode		
U1  a1 a2 b1 b2 cin Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ vinit_2bitpa		
U6  cin plot_v1		
U3  b2 plot_v1		
U2  b1 plot_v1		
U4  a2 plot_v1		
U5  a1 plot_v1		

.end
