* C:\Users\vinit\Desktop\SUMMATION-OF-COUNTER\1fullfinal\vinit_counter\vinit_counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/30/23 00:04:15

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ CLOCK Q00 vinit_dff		
U5  Net-_U5-Pad1_ CLOCK Q01 vinit_dff		
v1  clk GND pulse		
U3  clk CLOCK adc_bridge_1		
U4  clk plot_v1		
U6  q0 plot_v1		
U8  q1 plot_v1		
scmode1  SKY130mode		
X1  GND Q01 Q00 Net-_X1-Pad4_ Net-_U5-Pad1_ vinit_XOR		
v2  Net-_X1-Pad4_ GND 5		
U2  Q00 Q01 Net-_U13-Pad3_ Net-_U14-Pad3_ Net-_U2-Pad5_ S00 S01 S02 vinit_2bitpa		
U13  S00 CLOCK Net-_U13-Pad3_ vinit_dff		
U14  S01 CLOCK Net-_U14-Pad3_ vinit_dff		
U11  s0 plot_v1		
U10  s2 plot_v1		
U12  s1 plot_v1		
U15  Q00 Q01 S00 S01 S02 q0 q1 s0 s1 s2 dac_bridge_5		
X2  Net-_X1-Pad4_ Q00 GND Net-_U1-Pad1_ vinit_inverter		
U9  GND Net-_U2-Pad5_ adc_bridge_1		

.end
